
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package hash_array_pkg is

	type hash_array is array(integer range <>) of std_logic_vector(127 downto 0);

end hash_array_pkg;

package body hash_array_pkg is
 
end hash_array_pkg;